FILE_NAMING_RULE: %(entity_name)_entity.vhd
DESCRIPTION_START
This is the default template used for the creation of VHDL Entity files.
Template supplied by Mentor Graphics.
DESCRIPTION_END
-------------------------------------------------------------------------------
-- Title      : 
-- Project    : 
-------------------------------------------------------------------------------
-- File       : 
-- Author     : %(user)
-- Company    : Rohde & Schwarz
-- Last update: 
-- Platform   : PC
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date     Version     Author      Description
-------------------------------------------------------------------------------
%(entity)
