FILE_NAMING_RULE: %(class_name).svh
DESCRIPTION_START
This is the default template used for the creation of Class files.
Template supplied by Mentor Graphics.
DESCRIPTION_END
//
// Verilog class %(library).%(unit)
//
// Created:
//          by - %(user).%(group) (%(host))
//          at - %(time) %(date)
//
// using Mentor Graphics HDL Designer(TM) %(version)
//
%(classBody)
// ### Please start your Verilog code here ### 

endclass
