FILE_NAMING_RULE: %(entity_name)_%(arch_name).vhd
DESCRIPTION_START
This is the default template used for the creation of combined VHDL Architecture and Entity files.
Template supplied by Mentor Graphics.
DESCRIPTION_END
-------------------------------------------------------------------------------
-- Title      : 
-- Project    : 
-------------------------------------------------------------------------------
-- File       : %(entity_name)_%(arch_name).vhd
-- Author     : %(user)
-- Company    : Rohde & Schwarz
-- Last update: 
-- Platform   : PC
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date     Version     Author      Description
-------------------------------------------------------------------------------
%(entity)
--
%(architecture)
