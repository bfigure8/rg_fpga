-------------------------------------------------------------------------------
-- Title      : 
-- Project    : 
-------------------------------------------------------------------------------
-- File       : fpga_dac_a_rtl.vhd
-- Author     : steel_lake
-- Company    : DSO National Laboratories
-- Last update: 
-- Platform   : PC
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date     Version     Author      Description
-------------------------------------------------------------------------------
architecture rtl of fpga_dac_a is
begin
end architecture rtl;

