FILE_NAMING_RULE: %(program_name).sv
DESCRIPTION_START
This is the default template used for the creation of program files.
Template supplied by Mentor Graphics.
DESCRIPTION_END
//
// Verilog program %(library).%(unit)
//
// Created:
//          by - %(user).%(group) (%(host))
//          at - %(time) %(date)
//
// using Mentor Graphics HDL Designer(TM) %(version)
//
%(programBody)

// ### Please start your Verilog code here ### 
endprogram
