FILE_NAMING_RULE: %(interface_name).sv
DESCRIPTION_START
This is the default template used for the creation of Interface files.
Template supplied by Mentor Graphics.
DESCRIPTION_END
//
// Verilog interface %(library).%(unit)
//
// Created:
//          by - %(user).%(group) (%(host))
//          at - %(time) %(date)
//
// using Mentor Graphics HDL Designer(TM) %(version)
//
%(interfaceBody)

// ### Please start your Verilog code here ### 
endinterface
