FILE_NAMING_RULE: %(package_name).sv
DESCRIPTION_START
This is the default template used for the creation of Package files.
Template supplied by Mentor Graphics.
DESCRIPTION_END
//
// Verilog package %(library).%(unit)
//
// Created:
//          by - %(user).%(group) (%(host))
//          at - %(time) %(date)
//
// using Mentor Graphics HDL Designer(TM) %(version)
//
%(packageBody)
// ### Please start your Verilog code here ### 

endpackage
