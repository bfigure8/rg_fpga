FILE_NAMING_RULE: %(entity_name)_pkg_body.vhd
DESCRIPTION_START
This is the default template used for the creation of VHDL Package Body files.
Template supplied by Mentor Graphics.
DESCRIPTION_END
-------------------------------------------------------------------------------
-- Title      : 
-- Project    : 
-------------------------------------------------------------------------------
-- File       : 
-- Author     : %(user)
-- Company    : Rohde & Schwarz
-- Last update: 
-- Platform   : PC
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date     Version     Author      Description
-------------------------------------------------------------------------------
package body %(entity_name) is


end %(entity_name);