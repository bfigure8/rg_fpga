FILE_NAMING_RULE: %(module_name).v
DESCRIPTION_START
This is the default template used for the creation of Verilog Module files.
Template supplied by Mentor Graphics.
DESCRIPTION_END
//
// Verilog Module %(library).%(unit)
//
// Created:
//          by - %(user).%(group) (%(host))
//          at - %(time) %(date)
//
// using Mentor Graphics HDL Designer(TM) %(version)
//
%(moduleBody)
// ### Please start your Verilog code here ### 

endmodule
